*-----------------------------------------------------------------
* StrongARM sense latch for sharedDriveDiff feed
*-----------------------------------------------------------------
.subckt STRONGARM_INVERT sharedDriveP sharedDriveN comp_out vdd 0
.param COMP_WP=4u
.param COMP_WN=2u
.param COMP_L=0.13u
.param COMP_WP_CROSS={COMP_WP}
.param COMP_WN_TAIL={COMP_WN}
.param COMP_WN_LOAD={COMP_WN}
.param comp_l={COMP_L}
.param comp_wp_cross={COMP_WP_CROSS}
.param comp_wn_tail={COMP_WN_TAIL}
.param comp_wn_load={COMP_WN_LOAD}
Mpf1 comp_out sharedDriveP out_int vdd sky130_fd_pr__pfet_01v8__ss l={COMP_L} w={COMP_WP_CROSS} nf=1 ad={COMP_WP_CROSS*COMP_L} as={COMP_WP_CROSS*COMP_L} pd={2*(COMP_WP_CROSS+COMP_L)} ps={2*(COMP_WP_CROSS+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
Mpf2 comp_out sharedDriveN out_int vdd sky130_fd_pr__pfet_01v8__ss l={COMP_L} w={COMP_WP_CROSS} nf=1 ad={COMP_WP_CROSS*COMP_L} as={COMP_WP_CROSS*COMP_L} pd={2*(COMP_WP_CROSS+COMP_L)} ps={2*(COMP_WP_CROSS+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
Mpf3 out_int sharedDriveP mid vdd sky130_fd_pr__pfet_01v8__ss l={COMP_L} w={COMP_WP_CROSS} nf=1 ad={COMP_WP_CROSS*COMP_L} as={COMP_WP_CROSS*COMP_L} pd={2*(COMP_WP_CROSS+COMP_L)} ps={2*(COMP_WP_CROSS+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
Mpf4 out_int sharedDriveN mid vdd sky130_fd_pr__pfet_01v8__ss l={COMP_L} w={COMP_WP_CROSS} nf=1 ad={COMP_WP_CROSS*COMP_L} as={COMP_WP_CROSS*COMP_L} pd={2*(COMP_WP_CROSS+COMP_L)} ps={2*(COMP_WP_CROSS+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
Mnf1 comp_out mid 0 0 sky130_fd_pr__nfet_01v8__ss l={COMP_L} w={COMP_WN_TAIL} nf=1 ad={COMP_WN_TAIL*COMP_L} as={COMP_WN_TAIL*COMP_L} pd={2*(COMP_WN_TAIL+COMP_L)} ps={2*(COMP_WN_TAIL+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
Mnf2 comp_out comp_out 0 0 sky130_fd_pr__nfet_01v8__ss l={COMP_L} w={COMP_WN_LOAD} nf=1 ad={COMP_WN_LOAD*COMP_L} as={COMP_WN_LOAD*COMP_L} pd={2*(COMP_WN_LOAD+COMP_L)} ps={2*(COMP_WN_LOAD+COMP_L)} nrd=1 nrs=1 sa=0 sb=0 sd=0
.ends
